

package ALU_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"



`include "ALU_seqence_item.sv"
`include "sequence.sv"
`include "Sequencer.sv"
`include "Driver.sv"
`include "Monitor.sv"
`include "Agent.sv"
`include "Scoreborad.sv"
`include "Environment.sv"
`include "ALU_Test.sv"




endpackage


`include "interface.sv"